module and_gate(output o, input i1, i2, i3, i4);

assign o = i1 & i2 & i3 & i4;

endmodule
