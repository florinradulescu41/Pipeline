module imm_gen(input [31:0] in, output reg [31:0] out);

wire [9:0] sw; 

assign sw = {in[14:12], in[6:0]};

always @ (*) 
	begin
	case(sw)
		10'b0100000011: out <= {{21 {in[31]}}, in[30:25], in[24:21], in[20]};  
		10'b0000010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};  
		10'b1110010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};
		10'b1100010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};
		10'b1000010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};
		10'b0100010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};
		10'b0110010011: out <=  {{21 {in[31]}}, in[30:25], in[24:21], in[20]};
		10'b1010010011: out <=  {{21 {in[31]}}, in[30:25], in[11:8], in[7]};
		10'b0010010011: out <=  {{21 {in[31]}}, in[30:25], in[11:8], in[7]};
		10'b0100100011: out <=  {{21 {in[31]}}, in[30:25], in[11:8], in[7]};
		10'b0001100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
		10'b0011100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
		10'b1001100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
		10'b1011100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
		10'b1101100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
		10'b1111100011: out <=  {{20 {in[31]}}, in[7], in[30:25], in[11:8], 1'b0};
	endcase
	end

endmodule
