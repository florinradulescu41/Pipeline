module or_gate(output o, input i1, i2, i3, i4, i5, i6, i7, i8);

assign o = i1 | i2 | i3 | i4 | i5 | i6 | i7 | i8;

endmodule

