module not_gate(output o, input i);

assign o = ~ i;

endmodule
